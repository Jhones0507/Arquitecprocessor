library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity RegisterFile is
    Port ( 
				  Reset : in  STD_LOGIC;
				  rs1 : in  STD_LOGIC_VECTOR (5 downto 0);
				  rs2 : in  STD_LOGIC_VECTOR (5 downto 0);
				  rd : in  STD_LOGIC_VECTOR (5 downto 0);
				  DWR : in  STD_LOGIC_VECTOR (31 downto 0);
				  writeEnable : in  STD_LOGIC;
				  Crs1 : out  STD_LOGIC_VECTOR (31 downto 0);
				  Crs2 : out  STD_LOGIC_VECTOR (31 downto 0);
				  CRd : out  STD_LOGIC_VECTOR (31 downto 0)
			 );
end RegisterFile;

architecture Behavioral of RegisterFile is
type ram_type is array (0 to 39) of std_logic_vector (31 downto 0);
signal registro : ram_type := (
 "00000000000000000000000000000000","00000000000000000000000000000000",
 "00000000000000000000000000000000","00000000000000000000000000000000",
 "00000000000000000000000000000000","00000000000000000000000000000000",
 "00000000000000000000000000000000","00000000000000000000000000000000",
 "00000000000000000000000000000000","00000000000000000000000000000000",
 "00000000000000000000000000000000","00000000000000000000000000000000",
 "00000000000000000000000000000000","00000000000000000000000000000000",
 "00000000000000000000000000000000","00000000000000000000000000000000",
 "00000000000000000000000000000000","00000000000000000000000000000000",
 "00000000000000000000000000000000","00000000000000000000000000000000",
 "00000000000000000000000000000000","00000000000000000000000000000000",
 "00000000000000000000000000000000","00000000000000000000000000000000",
 "00000000000000000000000000000000","00000000000000000000000000000000",
 "00000000000000000000000000000000","00000000000000000000000000000000",
 "00000000000000000000000000000000","00000000000000000000000000000000",
 "00000000000000000000000000000000","00000000000000000000000000000000",
 "00000000000000000000000000000000","00000000000000000000000000000000",
 "00000000000000000000000000000000","00000000000000000000000000000000",
 "00000000000000000000000000000000","00000000000000000000000000000000",
 "00000000000000000000000000000000","00000000000000000000000000000000"
 ); 
begin

process(reset,rs1,rs2,rd,DWR,writeEnable)
 begin
 registro(0)<="00000000000000000000000000000000";
 if(Reset = '1')then
 Crs1 <= (others=>'0');
 Crs2 <= (others=>'0');
 CRd <= (others=>'0');
 registro <=(others => "00000000000000000000000000000000");
 else
 Crs1 <= registro(conv_integer(rs1));
 Crs2 <= registro(conv_integer(rs2));
 CRd <= registro(conv_integer(rd));
 if (writeEnable ='1' and rd/= "00000" )then
 registro(conv_integer(rd)) <= DWR ;
 end if;
 end if;
 end process;
end Behavioral;

